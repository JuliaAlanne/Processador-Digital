library verilog;
use verilog.vl_types.all;
entity altProcessor_vlg_vec_tst is
end altProcessor_vlg_vec_tst;
